//the difference between local and protected can be demonstrated in inheritance
